
//
// RISCV multi-cycle implementation.
//
// Module:      <module name>
//
// Description: <module description>
//
//

`include "rvm_constants.v"

module rvm_(

);



endmodule
