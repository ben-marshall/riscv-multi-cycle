
//
// RISCV multi-cycle implementation.
//
// Module:      axi_sram
//
// Description: A simple AXI SRAM module for testing.
//
//

`include "rvm_constants.v"

module axi_sram(

);



endmodule
